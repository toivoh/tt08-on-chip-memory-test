/*
 * Copyright (c) 2024 Toivo Henningsson
 * SPDX-License-Identifier: Apache-2.0
 */

`define ADDR_BITS 5
`define DATA_BITS 8
`define SERIAL_BITS 1
